magic
tech sky130A
magscale 1 2
timestamp 1729390267
<< obsli1 >>
rect 1104 2159 558808 349809
<< obsm1 >>
rect 934 2128 558808 349840
<< metal2 >>
rect 139950 0 140006 800
rect 419906 0 419962 800
<< obsm2 >>
rect 938 856 558698 349829
rect 938 800 139894 856
rect 140062 800 419850 856
rect 420018 800 558698 856
<< metal3 >>
rect 0 341640 800 341760
rect 559200 341640 560000 341760
rect 0 327224 800 327344
rect 559200 327224 560000 327344
rect 0 312808 800 312928
rect 559200 312808 560000 312928
rect 0 298392 800 298512
rect 559200 298392 560000 298512
rect 0 283976 800 284096
rect 559200 283976 560000 284096
rect 0 269560 800 269680
rect 559200 269560 560000 269680
rect 0 255144 800 255264
rect 559200 255144 560000 255264
rect 0 240728 800 240848
rect 559200 240728 560000 240848
rect 0 226312 800 226432
rect 559200 226312 560000 226432
rect 0 211896 800 212016
rect 559200 211896 560000 212016
rect 0 197480 800 197600
rect 559200 197480 560000 197600
rect 0 183064 800 183184
rect 559200 183064 560000 183184
rect 0 168648 800 168768
rect 559200 168648 560000 168768
rect 0 154232 800 154352
rect 559200 154232 560000 154352
rect 0 139816 800 139936
rect 559200 139816 560000 139936
rect 0 125400 800 125520
rect 559200 125400 560000 125520
rect 0 110984 800 111104
rect 559200 110984 560000 111104
rect 0 96568 800 96688
rect 559200 96568 560000 96688
rect 0 82152 800 82272
rect 559200 82152 560000 82272
rect 0 67736 800 67856
rect 559200 67736 560000 67856
rect 0 53320 800 53440
rect 559200 53320 560000 53440
rect 0 38904 800 39024
rect 559200 38904 560000 39024
rect 0 24488 800 24608
rect 559200 24488 560000 24608
rect 0 10072 800 10192
rect 559200 10072 560000 10192
<< obsm3 >>
rect 798 341840 559200 349825
rect 880 341560 559120 341840
rect 798 327424 559200 341560
rect 880 327144 559120 327424
rect 798 313008 559200 327144
rect 880 312728 559120 313008
rect 798 298592 559200 312728
rect 880 298312 559120 298592
rect 798 284176 559200 298312
rect 880 283896 559120 284176
rect 798 269760 559200 283896
rect 880 269480 559120 269760
rect 798 255344 559200 269480
rect 880 255064 559120 255344
rect 798 240928 559200 255064
rect 880 240648 559120 240928
rect 798 226512 559200 240648
rect 880 226232 559120 226512
rect 798 212096 559200 226232
rect 880 211816 559120 212096
rect 798 197680 559200 211816
rect 880 197400 559120 197680
rect 798 183264 559200 197400
rect 880 182984 559120 183264
rect 798 168848 559200 182984
rect 880 168568 559120 168848
rect 798 154432 559200 168568
rect 880 154152 559120 154432
rect 798 140016 559200 154152
rect 880 139736 559120 140016
rect 798 125600 559200 139736
rect 880 125320 559120 125600
rect 798 111184 559200 125320
rect 880 110904 559120 111184
rect 798 96768 559200 110904
rect 880 96488 559120 96768
rect 798 82352 559200 96488
rect 880 82072 559120 82352
rect 798 67936 559200 82072
rect 880 67656 559120 67936
rect 798 53520 559200 67656
rect 880 53240 559120 53520
rect 798 39104 559200 53240
rect 880 38824 559120 39104
rect 798 24688 559200 38824
rect 880 24408 559120 24688
rect 798 10272 559200 24408
rect 880 9992 559120 10272
rect 798 2143 559200 9992
<< metal4 >>
rect 4208 2128 4528 349840
rect 19568 2128 19888 349840
rect 34928 2128 35248 349840
rect 50288 2128 50608 349840
rect 65648 2128 65968 349840
rect 81008 2128 81328 349840
rect 96368 2128 96688 349840
rect 111728 2128 112048 349840
rect 127088 2128 127408 349840
rect 142448 2128 142768 349840
rect 157808 2128 158128 349840
rect 173168 2128 173488 349840
rect 188528 2128 188848 349840
rect 203888 2128 204208 349840
rect 219248 2128 219568 349840
rect 234608 2128 234928 349840
rect 249968 2128 250288 349840
rect 265328 2128 265648 349840
rect 280688 2128 281008 349840
rect 296048 2128 296368 349840
rect 311408 2128 311728 349840
rect 326768 2128 327088 349840
rect 342128 2128 342448 349840
rect 357488 2128 357808 349840
rect 372848 2128 373168 349840
rect 388208 2128 388528 349840
rect 403568 2128 403888 349840
rect 418928 2128 419248 349840
rect 434288 2128 434608 349840
rect 449648 2128 449968 349840
rect 465008 2128 465328 349840
rect 480368 2128 480688 349840
rect 495728 2128 496048 349840
rect 511088 2128 511408 349840
rect 526448 2128 526768 349840
rect 541808 2128 542128 349840
rect 557168 2128 557488 349840
<< labels >>
rlabel metal3 s 559200 10072 560000 10192 6 io_in[0]
port 1 nsew signal input
rlabel metal3 s 0 255144 800 255264 6 io_in[10]
port 2 nsew signal input
rlabel metal3 s 0 211896 800 212016 6 io_in[11]
port 3 nsew signal input
rlabel metal3 s 0 168648 800 168768 6 io_in[12]
port 4 nsew signal input
rlabel metal3 s 0 125400 800 125520 6 io_in[13]
port 5 nsew signal input
rlabel metal3 s 0 82152 800 82272 6 io_in[14]
port 6 nsew signal input
rlabel metal3 s 0 38904 800 39024 6 io_in[15]
port 7 nsew signal input
rlabel metal3 s 559200 53320 560000 53440 6 io_in[1]
port 8 nsew signal input
rlabel metal3 s 559200 96568 560000 96688 6 io_in[2]
port 9 nsew signal input
rlabel metal3 s 559200 139816 560000 139936 6 io_in[3]
port 10 nsew signal input
rlabel metal3 s 559200 183064 560000 183184 6 io_in[4]
port 11 nsew signal input
rlabel metal3 s 559200 226312 560000 226432 6 io_in[5]
port 12 nsew signal input
rlabel metal3 s 559200 269560 560000 269680 6 io_in[6]
port 13 nsew signal input
rlabel metal3 s 559200 312808 560000 312928 6 io_in[7]
port 14 nsew signal input
rlabel metal3 s 0 341640 800 341760 6 io_in[8]
port 15 nsew signal input
rlabel metal3 s 0 298392 800 298512 6 io_in[9]
port 16 nsew signal input
rlabel metal3 s 559200 38904 560000 39024 6 io_oeb[0]
port 17 nsew signal output
rlabel metal3 s 0 226312 800 226432 6 io_oeb[10]
port 18 nsew signal output
rlabel metal3 s 0 183064 800 183184 6 io_oeb[11]
port 19 nsew signal output
rlabel metal3 s 0 139816 800 139936 6 io_oeb[12]
port 20 nsew signal output
rlabel metal3 s 0 96568 800 96688 6 io_oeb[13]
port 21 nsew signal output
rlabel metal3 s 0 53320 800 53440 6 io_oeb[14]
port 22 nsew signal output
rlabel metal3 s 0 10072 800 10192 6 io_oeb[15]
port 23 nsew signal output
rlabel metal3 s 559200 82152 560000 82272 6 io_oeb[1]
port 24 nsew signal output
rlabel metal3 s 559200 125400 560000 125520 6 io_oeb[2]
port 25 nsew signal output
rlabel metal3 s 559200 168648 560000 168768 6 io_oeb[3]
port 26 nsew signal output
rlabel metal3 s 559200 211896 560000 212016 6 io_oeb[4]
port 27 nsew signal output
rlabel metal3 s 559200 255144 560000 255264 6 io_oeb[5]
port 28 nsew signal output
rlabel metal3 s 559200 298392 560000 298512 6 io_oeb[6]
port 29 nsew signal output
rlabel metal3 s 559200 341640 560000 341760 6 io_oeb[7]
port 30 nsew signal output
rlabel metal3 s 0 312808 800 312928 6 io_oeb[8]
port 31 nsew signal output
rlabel metal3 s 0 269560 800 269680 6 io_oeb[9]
port 32 nsew signal output
rlabel metal3 s 559200 24488 560000 24608 6 io_out[0]
port 33 nsew signal output
rlabel metal3 s 0 240728 800 240848 6 io_out[10]
port 34 nsew signal output
rlabel metal3 s 0 197480 800 197600 6 io_out[11]
port 35 nsew signal output
rlabel metal3 s 0 154232 800 154352 6 io_out[12]
port 36 nsew signal output
rlabel metal3 s 0 110984 800 111104 6 io_out[13]
port 37 nsew signal output
rlabel metal3 s 0 67736 800 67856 6 io_out[14]
port 38 nsew signal output
rlabel metal3 s 0 24488 800 24608 6 io_out[15]
port 39 nsew signal output
rlabel metal3 s 559200 67736 560000 67856 6 io_out[1]
port 40 nsew signal output
rlabel metal3 s 559200 110984 560000 111104 6 io_out[2]
port 41 nsew signal output
rlabel metal3 s 559200 154232 560000 154352 6 io_out[3]
port 42 nsew signal output
rlabel metal3 s 559200 197480 560000 197600 6 io_out[4]
port 43 nsew signal output
rlabel metal3 s 559200 240728 560000 240848 6 io_out[5]
port 44 nsew signal output
rlabel metal3 s 559200 283976 560000 284096 6 io_out[6]
port 45 nsew signal output
rlabel metal3 s 559200 327224 560000 327344 6 io_out[7]
port 46 nsew signal output
rlabel metal3 s 0 327224 800 327344 6 io_out[8]
port 47 nsew signal output
rlabel metal3 s 0 283976 800 284096 6 io_out[9]
port 48 nsew signal output
rlabel metal4 s 4208 2128 4528 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 127088 2128 127408 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 157808 2128 158128 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 188528 2128 188848 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 219248 2128 219568 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 249968 2128 250288 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 280688 2128 281008 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 311408 2128 311728 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 342128 2128 342448 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 372848 2128 373168 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 403568 2128 403888 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 434288 2128 434608 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 465008 2128 465328 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 495728 2128 496048 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 526448 2128 526768 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 557168 2128 557488 349840 6 vccd1
port 49 nsew power bidirectional
rlabel metal4 s 19568 2128 19888 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 142448 2128 142768 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 173168 2128 173488 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 203888 2128 204208 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 234608 2128 234928 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 265328 2128 265648 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 296048 2128 296368 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 326768 2128 327088 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 357488 2128 357808 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 388208 2128 388528 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 418928 2128 419248 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 449648 2128 449968 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 480368 2128 480688 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 511088 2128 511408 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal4 s 541808 2128 542128 349840 6 vssd1
port 50 nsew ground bidirectional
rlabel metal2 s 139950 0 140006 800 6 wb_clk_i
port 51 nsew signal input
rlabel metal2 s 419906 0 419962 800 6 wb_rst_i
port 52 nsew signal input
<< properties >>
string FIXED_BBOX 0 0 560000 352000
string LEFclass BLOCK
string LEFview TRUE
string GDS_END 52161560
string GDS_FILE /home/ngk/unic_cass_ic/uniccass_example/openlane/user_proj_example/runs/24_10_20_07_32/results/signoff/user_proj_example.magic.gds
string GDS_START 341820
<< end >>

